
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.uft_pkg.all;

entity entity_name is
    --generic (
    --    GEN1 : natural := 42042;
    --);
    port (
        -- clk and reset
        ------------------------------------------------------------------------
        clk     : in    std_logic;
        rst_n   : in    std_logic

    );
end entity entity_name;

architecture structural of entity_name is

begin

end architecture structural;